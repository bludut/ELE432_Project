
module Pll_50_to_25 (
	clk_clk,
	reset_reset_n,
	pll_0_outclk0_clk);	

	input		clk_clk;
	input		reset_reset_n;
	output		pll_0_outclk0_clk;
endmodule
