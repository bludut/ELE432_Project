library IEEE;
use IEEE.std_logic_1164.All;
use IEEE.numeric_std.All;
use IEEE.std_logic_unsigned.All;
entity Wall_Cars_Generator is
	Generic(
				g_Total_Row : integer := 480;
				g_Total_Column : integer := 640
				);
	Port(
			i_Dist_Ena : in Std_logic;
			i_Row_Num : in std_logic_vector (9 downto 0) ;
			i_Column_Num : in std_logic_vector (9 downto 0);
			i_Pos_X : in std_logic_vector(9 downto 0);
			i_Pos_Y : in std_logic_vector(9 downto 0);
			
			Cnst_2Car : in std_logic_vector(9 downto 0);
			Cnst_3Car : in std_logic_vector(9 downto 0);
			Cnst_4Car : in std_logic_vector(9 downto 0);		
			
			o_Red : out std_logic_vector (7 downto 0);
			o_Green : out std_logic_vector (7 downto 0);
			o_Blue : out std_logic_vector (7 downto 0);
			o_Disp_Ena : out std_logic
			);
end Wall_Cars_Generator;


architecture arch of Wall_Cars_Generator is

	------------------------------------------------------------------
	-- WALL GENERATOR
	------------------------------------------------------------------
	component Wall_Generator is
	Generic(
				g_Total_Row : integer := 480;
				g_Total_Column : integer := 640
				);
	Port(
			i_Dist_Ena : in Std_logic;
			i_Row_Num : in std_logic_vector (9 downto 0) ;
			i_Column_Num : in std_logic_vector (9 downto 0);
			i_Pos_X : in std_logic_vector(9 downto 0);
			i_Pos_Y : in std_logic_vector(9 downto 0);
			
			o_Red : out std_logic_vector (7 downto 0);
			o_Green : out std_logic_vector (7 downto 0);
			o_Blue : out std_logic_vector (7 downto 0);
			o_Disp_Ena : out std_logic
			);
	end component Wall_Generator;
		
--	constant Cnst_2Car : std_logic_vector(9 downto 0) := "00" & X"C8";		-- Second Car offset = 200 
--	constant Cnst_3Car : std_logic_vector(9 downto 0) := "00" & X"C8";		-- Second Car offset = 200
--	constant Cnst_3Car : std_logic_vector(9 downto 0) := "00" & X"C8";		-- Second Car offset = 200

	

	signal o_Car_Disp_Ena : std_logic_vector(3 downto 0);
begin

	-- First Car
Car1:component Wall_Generator 
	Generic map(
				g_Total_Row => 480,
				g_Total_Column => 640
				)
	Port map(
			i_Dist_Ena => i_Dist_Ena,
			i_Row_Num => i_Row_Num,
			i_Column_Num => i_Column_Num,
			i_Pos_X => i_Pos_X,
			i_Pos_Y => i_Pos_Y,
			
			o_Red => o_Red,
			o_Green => o_Green,
			o_Blue => o_Blue,
			o_Disp_Ena => o_Car_Disp_Ena(0)
			);
			
	-- Second Car
Car2:component Wall_Generator 
	Generic map(
				g_Total_Row => 480,
				g_Total_Column => 640
				)
	Port map(
			i_Dist_Ena => i_Dist_Ena,
			i_Row_Num => i_Row_Num,
			i_Column_Num => i_Column_Num,
			i_Pos_X => i_Pos_X,
			i_Pos_Y => i_Pos_Y + Cnst_2Car,
			
			o_Red => open,
			o_Green => open,
			o_Blue => open,
			o_Disp_Ena => o_Car_Disp_Ena(1)
			);
			
	-- Third Car
Car3:component Wall_Generator 
	Generic map(
				g_Total_Row => 480,
				g_Total_Column => 640
				)
	Port map(
			i_Dist_Ena => i_Dist_Ena,
			i_Row_Num => i_Row_Num,
			i_Column_Num => i_Column_Num,
			i_Pos_X => i_Pos_X,
			i_Pos_Y => i_Pos_Y + Cnst_3Car,
			
			o_Red => open,
			o_Green => open,
			o_Blue => open,
			o_Disp_Ena => o_Car_Disp_Ena(2)
			);
			
	-- 4th Car
Car4:component Wall_Generator 
	Generic map(
				g_Total_Row => 480,
				g_Total_Column => 640
				)
	Port map(
			i_Dist_Ena => i_Dist_Ena,
			i_Row_Num => i_Row_Num,
			i_Column_Num => i_Column_Num,
			i_Pos_X => i_Pos_X,	
			i_Pos_Y => i_Pos_Y + Cnst_4Car,
			
			o_Red => open,
			o_Green => open,
			o_Blue => open,
			o_Disp_Ena => o_Car_Disp_Ena(3)
			);
			
			
-- OR'ed display enable
	o_Disp_Ena <=  o_Car_Disp_Ena(0) or
						o_Car_Disp_Ena(1) or
						o_Car_Disp_Ena(2) or
						o_Car_Disp_Ena(3);
				

end arch;